library	ieee;
use	ieee.std_logic_1164.all;
use	ieee.numeric_std.all;

package	mips_pkg	is
	-- Declaracao	de	componentes
	component breg_ula is
		generic	(	WSIZE	:	natural	:=	32);
		port(
			rs,rt, rd : in std_logic_vector(4 downto 0);
			we, clk : in std_logic;
			din : in std_logic_vector(31 downto 0);
			func : in std_logic_vector(5 downto 0);
			opula : in std_logic_vector(1 downto 0);
			dout  : out std_logic_vector(31 downto 0);
			zero : out std_logic
		);
	end component;
	
	component	ula	is
		generic	(	WSIZE	:	natural	:=	32);
		port	(	
			ulop :	in	std_logic_vector(3	downto	0);
			A,	B :	in	std_logic_vector(WSIZE-1	downto	0);	
			aluout:	out	std_logic_vector(WSIZE-1	downto	0);	
			zero :	out	std_logic	
			);
	end	component;
	
	component	c_ula	is
		port	(
			func	 :	in	std_logic_vector(5	downto	0);
			opUla :	in	std_logic_vector(1	downto	0);
			ctrula	 :	out	std_logic_vector(3	downto	0)
			);
	end	component;
	
	component	breg	is
		generic	(	WSIZE	:	natural	:=	32;
			ISIZE	:	natural	:=	5;
			BREGSIZE	:	natural	:=	32	);
		port	
			(
			clk :	in		std_logic;
			we :	in		std_logic;
			rs :	in		std_logic_vector(ISIZE-1	downto	0);
			rt :	in		std_logic_vector(ISIZE-1	downto	0);
			rd :	in		std_logic_vector(ISIZE-1	downto	0);
			d_in :	in		std_logic_vector(WSIZE-1	downto	0);
			regA	 :	out	std_logic_vector(WSIZE-1	downto	0);
			regB	 :	out	std_logic_vector(WSIZE-1	downto	0)
			);
	end	component;
	
	component somador is 
		generic	(	WSIZE	:	natural	:=	32);
		port(
			clk : in std_logic;
			A, B : in std_logic_vector ((WSIZE - 1) downto 0);

			result : out std_logic_vector ((WSIZE - 1) downto 0)
		);
	end component;
	
	component pc is
		generic	(	WSIZE	:	natural	:=	32);
		port(
			clk : in std_logic;
			input : in std_logic_vector ((WSIZE - 1) downto 0);

			output : out std_logic_vesctor (7 downto 0)
		);
	end component;
	
	component multiplexador_5_bits is
		port(
			selector : in std_logic;
			opt0, opt1 : in std_logic_vector (4 downto 0);
			result : out std_logic_vector (4 downto 0)
		);
	end component;

	component memory_instruction is
		port(
			address	: in std_logic_vector(7 downto 0);
			clock		: in std_logic;
			q		   : out std_logic_vector(31 downto 0)
		);
	end component;

	component control is
		port(
			opcode : in std_logic_vector(5 downto 0),
			RegDst : out std_logic;
			Jump : out std_logic;
			Brench : out std_logic;
			MemRead : out std_logic;
			MemtoReg : out std_logic;
			MemWrite : out std_logic;
			ALUOp : out std_logic_vector(1 downto 0);
			ALUSrc : out std_logic
		);
	end component;
	
	component data_memory is
		port(
			address	: in std_logic_vector(7 downto 0);
			clock		: in std_logic;
			data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			wren		: IN STD_LOGIC ;
			q		   : out std_logic_vector(31 downto 0)
		);
	end component;
	
	-- Controle	ULAmips
	constant	ULA_AND :	std_logic_vector(3	downto	0)	:=	"0000";	-- 0
	constant	ULA_OR :	std_logic_vector(3	downto	0)	:=	"0001";	-- 1
	constant	ULA_ADD :	std_logic_vector(3	downto	0)	:=	"0010";	-- 2
	constant	ULA_SUB :	std_logic_vector(3	downto	0)	:=	"0110";	-- 6
	constant	ULA_SLT :	std_logic_vector(3	downto	0)	:=	"0111";	-- 7
	constant	ULA_NOR :	std_logic_vector(3	downto	0)	:=	"1100";	-- 12
	constant	ULA_UKW :	std_logic_vector(3	downto	0)	:=	"XXXX";
end	mips_pkg;